module GC_Read ( input clk , input POLL , input GC_enable , input wire button2 ,
    output reg [15:0] GCBD , output reg GCpollend = 0 , output reg connected = 0 , output reg [2:0] connection_type = 3'b000 ,
    output reg [15:0] GCLA , output reg [15:0] GCRA , output reg [15:0] GCTA
);                                                                                      
reg prev_POLL = 1; reg [9:0] count = 0;  reg NSOCal = 0;
reg [6:0] bit_count = 7'd82;
reg signed [8:0] offsetx = 0; reg signed [8:0] offsety = 0; reg signed [8:0] offsetcx = 0; reg signed [8:0] offsetcy = 0; reg [8:0] offsetLT = 0; reg [8:0] offsetRT = 0;
reg signed [8:0] xcal = 0; reg signed [8:0] ycal = 0; reg signed [8:0] cxcal = 0; reg signed [8:0] cycal = 0;
reg [7:0] x; reg [7:0] y; reg [7:0] cx; reg [7:0] cy; reg [7:0] LAT; reg [7:0] RAT; 
always @ ( posedge clk ) begin //scale the output, using an approximation
    
    xcal  <= $signed({1'b0,GCdata[48:41]})-$signed(offsetx);
    ycal  <= $signed({1'b0,GCdata[40:33]})-$signed(offsety);
    cxcal <= $signed({1'b0,GCdata[32:25]})-$signed(offsetcx);
    cycal <= $signed({1'b0,GCdata[24:17]})-$signed(offsetcy);

case ( xcal )8'd0: x <= 8'd33;8'd1: x <= 8'd34;8'd2: x <= 8'd34;8'd3: x <= 8'd35;8'd4: x <= 8'd36;8'd5: x <= 8'd37;8'd6: x <= 8'd37;8'd7: x <= 8'd38;8'd8: x <= 8'd39;8'd9: x <= 8'd40;8'd10: x <= 8'd40;8'd11: x <= 8'd41;8'd12: x <= 8'd42;8'd13: x <= 8'd43;8'd14: x <= 8'd43;8'd15: x <= 8'd44;8'd16: x <= 8'd45;8'd17: x <= 8'd46;8'd18: x <= 8'd46;8'd19: x <= 8'd47;8'd20: x <= 8'd48;8'd21: x <= 8'd49;8'd22: x <= 8'd49;8'd23: x <= 8'd50;8'd24: x <= 8'd51;8'd25: x <= 8'd52;8'd26: x <= 8'd52;8'd27: x <= 8'd53;8'd28: x <= 8'd54;8'd29: x <= 8'd54;8'd30: x <= 8'd55;8'd31: x <= 8'd56;8'd32: x <= 8'd57;8'd33: x <= 8'd57;8'd34: x <= 8'd58;8'd35: x <= 8'd59;8'd36: x <= 8'd60;8'd37: x <= 8'd60;8'd38: x <= 8'd61;8'd39: x <= 8'd62;8'd40: x <= 8'd63;8'd41: x <= 8'd63;8'd42: x <= 8'd64;8'd43: x <= 8'd65;8'd44: x <= 8'd66;8'd45: x <= 8'd66;8'd46: x <= 8'd67;8'd47: x <= 8'd68;8'd48: x <= 8'd69;8'd49: x <= 8'd69;8'd50: x <= 8'd70;8'd51: x <= 8'd71;8'd52: x <= 8'd71;8'd53: x <= 8'd72;8'd54: x <= 8'd73;8'd55: x <= 8'd74;8'd56: x <= 8'd74;8'd57: x <= 8'd75;8'd58: x <= 8'd76;8'd59: x <= 8'd77;8'd60: x <= 8'd77;8'd61: x <= 8'd78;8'd62: x <= 8'd79;8'd63: x <= 8'd80;8'd64: x <= 8'd80;8'd65: x <= 8'd81;8'd66: x <= 8'd82;8'd67: x <= 8'd83;8'd68: x <= 8'd83;8'd69: x <= 8'd84;8'd70: x <= 8'd85;8'd71: x <= 8'd86;8'd72: x <= 8'd86;8'd73: x <= 8'd87;8'd74: x <= 8'd88;8'd75: x <= 8'd89;8'd76: x <= 8'd89;8'd77: x <= 8'd90;8'd78: x <= 8'd91;8'd79: x <= 8'd91;8'd80: x <= 8'd92;8'd81: x <= 8'd93;8'd82: x <= 8'd94;8'd83: x <= 8'd94;8'd84: x <= 8'd95;8'd85: x <= 8'd96;8'd86: x <= 8'd97;8'd87: x <= 8'd97;8'd88: x <= 8'd98;8'd89: x <= 8'd99;8'd90: x <= 8'd100;8'd91: x <= 8'd100;8'd92: x <= 8'd101;8'd93: x <= 8'd102;8'd94: x <= 8'd103;8'd95: x <= 8'd103;8'd96: x <= 8'd104;8'd97: x <= 8'd105;8'd98: x <= 8'd106;8'd99: x <= 8'd106;8'd100: x <= 8'd107;8'd101: x <= 8'd108;8'd102: x <= 8'd108;8'd103: x <= 8'd109;8'd104: x <= 8'd110;8'd105: x <= 8'd111;8'd106: x <= 8'd111;8'd107: x <= 8'd112;8'd108: x <= 8'd113;8'd109: x <= 8'd114;8'd110: x <= 8'd114;8'd111: x <= 8'd115;8'd112: x <= 8'd116;8'd113: x <= 8'd117;8'd114: x <= 8'd117;8'd115: x <= 8'd118;8'd116: x <= 8'd119;8'd117: x <= 8'd120;8'd118: x <= 8'd120;8'd119: x <= 8'd121;8'd120: x <= 8'd122;8'd121: x <= 8'd123;8'd122: x <= 8'd123;8'd123: x <= 8'd124;8'd124: x <= 8'd125;8'd125: x <= 8'd126;8'd126: x <= 8'd126;8'd127: x <= 8'd127;8'd128: x <= 8'd128;8'd129: x <= 8'd128;8'd130: x <= 8'd129;8'd131: x <= 8'd130;8'd132: x <= 8'd131;8'd133: x <= 8'd131;8'd134: x <= 8'd132;8'd135: x <= 8'd133;8'd136: x <= 8'd134;8'd137: x <= 8'd134;8'd138: x <= 8'd135;8'd139: x <= 8'd136;8'd140: x <= 8'd137;8'd141: x <= 8'd137;8'd142: x <= 8'd138;8'd143: x <= 8'd139;8'd144: x <= 8'd140;8'd145: x <= 8'd140;8'd146: x <= 8'd141;8'd147: x <= 8'd142;8'd148: x <= 8'd143;8'd149: x <= 8'd143;8'd150: x <= 8'd144;8'd151: x <= 8'd145;8'd152: x <= 8'd146;8'd153: x <= 8'd146;8'd154: x <= 8'd147;8'd155: x <= 8'd148;8'd156: x <= 8'd148;8'd157: x <= 8'd149;8'd158: x <= 8'd150;8'd159: x <= 8'd151;8'd160: x <= 8'd151;8'd161: x <= 8'd152;8'd162: x <= 8'd153;8'd163: x <= 8'd154;8'd164: x <= 8'd154;8'd165: x <= 8'd155;8'd166: x <= 8'd156;8'd167: x <= 8'd157;8'd168: x <= 8'd157;8'd169: x <= 8'd158;8'd170: x <= 8'd159;8'd171: x <= 8'd160;8'd172: x <= 8'd160;8'd173: x <= 8'd161;8'd174: x <= 8'd162;8'd175: x <= 8'd163;8'd176: x <= 8'd163;8'd177: x <= 8'd164;8'd178: x <= 8'd165;8'd179: x <= 8'd165;8'd180: x <= 8'd166;8'd181: x <= 8'd167;8'd182: x <= 8'd168;8'd183: x <= 8'd168;8'd184: x <= 8'd169;8'd185: x <= 8'd170;8'd186: x <= 8'd171;8'd187: x <= 8'd171;8'd188: x <= 8'd172;8'd189: x <= 8'd173;8'd190: x <= 8'd174;8'd191: x <= 8'd174;8'd192: x <= 8'd175;8'd193: x <= 8'd176;8'd194: x <= 8'd177;8'd195: x <= 8'd177;8'd196: x <= 8'd178;8'd197: x <= 8'd179;8'd198: x <= 8'd180;8'd199: x <= 8'd180;8'd200: x <= 8'd181;8'd201: x <= 8'd182;8'd202: x <= 8'd183;8'd203: x <= 8'd183;8'd204: x <= 8'd184;8'd205: x <= 8'd185;8'd206: x <= 8'd185;8'd207: x <= 8'd186;8'd208: x <= 8'd187;8'd209: x <= 8'd188;8'd210: x <= 8'd188;8'd211: x <= 8'd189;8'd212: x <= 8'd190;8'd213: x <= 8'd191;8'd214: x <= 8'd191;8'd215: x <= 8'd192;8'd216: x <= 8'd193;8'd217: x <= 8'd194;8'd218: x <= 8'd194;8'd219: x <= 8'd195;8'd220: x <= 8'd196;8'd221: x <= 8'd197;8'd222: x <= 8'd197;8'd223: x <= 8'd198;8'd224: x <= 8'd199;8'd225: x <= 8'd200;8'd226: x <= 8'd200;8'd227: x <= 8'd201;8'd228: x <= 8'd202;8'd229: x <= 8'd202;8'd230: x <= 8'd203;8'd231: x <= 8'd204;8'd232: x <= 8'd205;8'd233: x <= 8'd205;8'd234: x <= 8'd206;8'd235: x <= 8'd207;8'd236: x <= 8'd208;8'd237: x <= 8'd208;8'd238: x <= 8'd209;8'd239: x <= 8'd210;8'd240: x <= 8'd211;8'd241: x <= 8'd211;8'd242: x <= 8'd212;8'd243: x <= 8'd213;8'd244: x <= 8'd214;8'd245: x <= 8'd214;8'd246: x <= 8'd215;8'd247: x <= 8'd216;8'd248: x <= 8'd217;8'd249: x <= 8'd217;8'd250: x <= 8'd218;8'd251: x <= 8'd219;8'd252: x <= 8'd220;8'd253: x <= 8'd220;8'd254: x <= 8'd221;8'd255: x <= 8'd222;default: x<=8'd127; endcase case ( ycal )8'd0: y <= 8'd33;8'd1: y <= 8'd34;8'd2: y <= 8'd34;8'd3: y <= 8'd35;8'd4: y <= 8'd36;8'd5: y <= 8'd37;8'd6: y <= 8'd37;8'd7: y <= 8'd38;8'd8: y <= 8'd39;8'd9: y <= 8'd40;8'd10: y <= 8'd40;8'd11: y <= 8'd41;8'd12: y <= 8'd42;8'd13: y <= 8'd43;8'd14: y <= 8'd43;8'd15: y <= 8'd44;8'd16: y <= 8'd45;8'd17: y <= 8'd46;8'd18: y <= 8'd46;8'd19: y <= 8'd47;8'd20: y <= 8'd48;8'd21: y <= 8'd49;8'd22: y <= 8'd49;8'd23: y <= 8'd50;8'd24: y <= 8'd51;8'd25: y <= 8'd52;8'd26: y <= 8'd52;8'd27: y <= 8'd53;8'd28: y <= 8'd54;8'd29: y <= 8'd54;8'd30: y <= 8'd55;8'd31: y <= 8'd56;8'd32: y <= 8'd57;8'd33: y <= 8'd57;8'd34: y <= 8'd58;8'd35: y <= 8'd59;8'd36: y <= 8'd60;8'd37: y <= 8'd60;8'd38: y <= 8'd61;8'd39: y <= 8'd62;8'd40: y <= 8'd63;8'd41: y <= 8'd63;8'd42: y <= 8'd64;8'd43: y <= 8'd65;8'd44: y <= 8'd66;8'd45: y <= 8'd66;8'd46: y <= 8'd67;8'd47: y <= 8'd68;8'd48: y <= 8'd69;8'd49: y <= 8'd69;8'd50: y <= 8'd70;8'd51: y <= 8'd71;8'd52: y <= 8'd71;8'd53: y <= 8'd72;8'd54: y <= 8'd73;8'd55: y <= 8'd74;8'd56: y <= 8'd74;8'd57: y <= 8'd75;8'd58: y <= 8'd76;8'd59: y <= 8'd77;8'd60: y <= 8'd77;8'd61: y <= 8'd78;8'd62: y <= 8'd79;8'd63: y <= 8'd80;8'd64: y <= 8'd80;8'd65: y <= 8'd81;8'd66: y <= 8'd82;8'd67: y <= 8'd83;8'd68: y <= 8'd83;8'd69: y <= 8'd84;8'd70: y <= 8'd85;8'd71: y <= 8'd86;8'd72: y <= 8'd86;8'd73: y <= 8'd87;8'd74: y <= 8'd88;8'd75: y <= 8'd89;8'd76: y <= 8'd89;8'd77: y <= 8'd90;8'd78: y <= 8'd91;8'd79: y <= 8'd91;8'd80: y <= 8'd92;8'd81: y <= 8'd93;8'd82: y <= 8'd94;8'd83: y <= 8'd94;8'd84: y <= 8'd95;8'd85: y <= 8'd96;8'd86: y <= 8'd97;8'd87: y <= 8'd97;8'd88: y <= 8'd98;8'd89: y <= 8'd99;8'd90: y <= 8'd100;8'd91: y <= 8'd100;8'd92: y <= 8'd101;8'd93: y <= 8'd102;8'd94: y <= 8'd103;8'd95: y <= 8'd103;8'd96: y <= 8'd104;8'd97: y <= 8'd105;8'd98: y <= 8'd106;8'd99: y <= 8'd106;8'd100: y <= 8'd107;8'd101: y <= 8'd108;8'd102: y <= 8'd108;8'd103: y <= 8'd109;8'd104: y <= 8'd110;8'd105: y <= 8'd111;8'd106: y <= 8'd111;8'd107: y <= 8'd112;8'd108: y <= 8'd113;8'd109: y <= 8'd114;8'd110: y <= 8'd114;8'd111: y <= 8'd115;8'd112: y <= 8'd116;8'd113: y <= 8'd117;8'd114: y <= 8'd117;8'd115: y <= 8'd118;8'd116: y <= 8'd119;8'd117: y <= 8'd120;8'd118: y <= 8'd120;8'd119: y <= 8'd121;8'd120: y <= 8'd122;8'd121: y <= 8'd123;8'd122: y <= 8'd123;8'd123: y <= 8'd124;8'd124: y <= 8'd125;8'd125: y <= 8'd126;8'd126: y <= 8'd126;8'd127: y <= 8'd127;8'd128: y <= 8'd128;8'd129: y <= 8'd128;8'd130: y <= 8'd129;8'd131: y <= 8'd130;8'd132: y <= 8'd131;8'd133: y <= 8'd131;8'd134: y <= 8'd132;8'd135: y <= 8'd133;8'd136: y <= 8'd134;8'd137: y <= 8'd134;8'd138: y <= 8'd135;8'd139: y <= 8'd136;8'd140: y <= 8'd137;8'd141: y <= 8'd137;8'd142: y <= 8'd138;8'd143: y <= 8'd139;8'd144: y <= 8'd140;8'd145: y <= 8'd140;8'd146: y <= 8'd141;8'd147: y <= 8'd142;8'd148: y <= 8'd143;8'd149: y <= 8'd143;8'd150: y <= 8'd144;8'd151: y <= 8'd145;8'd152: y <= 8'd146;8'd153: y <= 8'd146;8'd154: y <= 8'd147;8'd155: y <= 8'd148;8'd156: y <= 8'd148;8'd157: y <= 8'd149;8'd158: y <= 8'd150;8'd159: y <= 8'd151;8'd160: y <= 8'd151;8'd161: y <= 8'd152;8'd162: y <= 8'd153;8'd163: y <= 8'd154;8'd164: y <= 8'd154;8'd165: y <= 8'd155;8'd166: y <= 8'd156;8'd167: y <= 8'd157;8'd168: y <= 8'd157;8'd169: y <= 8'd158;8'd170: y <= 8'd159;8'd171: y <= 8'd160;8'd172: y <= 8'd160;8'd173: y <= 8'd161;8'd174: y <= 8'd162;8'd175: y <= 8'd163;8'd176: y <= 8'd163;8'd177: y <= 8'd164;8'd178: y <= 8'd165;8'd179: y <= 8'd165;8'd180: y <= 8'd166;8'd181: y <= 8'd167;8'd182: y <= 8'd168;8'd183: y <= 8'd168;8'd184: y <= 8'd169;8'd185: y <= 8'd170;8'd186: y <= 8'd171;8'd187: y <= 8'd171;8'd188: y <= 8'd172;8'd189: y <= 8'd173;8'd190: y <= 8'd174;8'd191: y <= 8'd174;8'd192: y <= 8'd175;8'd193: y <= 8'd176;8'd194: y <= 8'd177;8'd195: y <= 8'd177;8'd196: y <= 8'd178;8'd197: y <= 8'd179;8'd198: y <= 8'd180;8'd199: y <= 8'd180;8'd200: y <= 8'd181;8'd201: y <= 8'd182;8'd202: y <= 8'd183;8'd203: y <= 8'd183;8'd204: y <= 8'd184;8'd205: y <= 8'd185;8'd206: y <= 8'd185;8'd207: y <= 8'd186;8'd208: y <= 8'd187;8'd209: y <= 8'd188;8'd210: y <= 8'd188;8'd211: y <= 8'd189;8'd212: y <= 8'd190;8'd213: y <= 8'd191;8'd214: y <= 8'd191;8'd215: y <= 8'd192;8'd216: y <= 8'd193;8'd217: y <= 8'd194;8'd218: y <= 8'd194;8'd219: y <= 8'd195;8'd220: y <= 8'd196;8'd221: y <= 8'd197;8'd222: y <= 8'd197;8'd223: y <= 8'd198;8'd224: y <= 8'd199;8'd225: y <= 8'd200;8'd226: y <= 8'd200;8'd227: y <= 8'd201;8'd228: y <= 8'd202;8'd229: y <= 8'd202;8'd230: y <= 8'd203;8'd231: y <= 8'd204;8'd232: y <= 8'd205;8'd233: y <= 8'd205;8'd234: y <= 8'd206;8'd235: y <= 8'd207;8'd236: y <= 8'd208;8'd237: y <= 8'd208;8'd238: y <= 8'd209;8'd239: y <= 8'd210;8'd240: y <= 8'd211;8'd241: y <= 8'd211;8'd242: y <= 8'd212;8'd243: y <= 8'd213;8'd244: y <= 8'd214;8'd245: y <= 8'd214;8'd246: y <= 8'd215;8'd247: y <= 8'd216;8'd248: y <= 8'd217;8'd249: y <= 8'd217;8'd250: y <= 8'd218;8'd251: y <= 8'd219;8'd252: y <= 8'd220;8'd253: y <= 8'd220;8'd254: y <= 8'd221;8'd255: y <= 8'd222;default: y<=8'd127; endcase case ( cxcal )8'd0: cx <= 8'd33;8'd1: cx <= 8'd34;8'd2: cx <= 8'd34;8'd3: cx <= 8'd35;8'd4: cx <= 8'd36;8'd5: cx <= 8'd37;8'd6: cx <= 8'd37;8'd7: cx <= 8'd38;8'd8: cx <= 8'd39;8'd9: cx <= 8'd40;8'd10: cx <= 8'd40;8'd11: cx <= 8'd41;8'd12: cx <= 8'd42;8'd13: cx <= 8'd43;8'd14: cx <= 8'd43;8'd15: cx <= 8'd44;8'd16: cx <= 8'd45;8'd17: cx <= 8'd46;8'd18: cx <= 8'd46;8'd19: cx <= 8'd47;8'd20: cx <= 8'd48;8'd21: cx <= 8'd49;8'd22: cx <= 8'd49;8'd23: cx <= 8'd50;8'd24: cx <= 8'd51;8'd25: cx <= 8'd52;8'd26: cx <= 8'd52;8'd27: cx <= 8'd53;8'd28: cx <= 8'd54;8'd29: cx <= 8'd54;8'd30: cx <= 8'd55;8'd31: cx <= 8'd56;8'd32: cx <= 8'd57;8'd33: cx <= 8'd57;8'd34: cx <= 8'd58;8'd35: cx <= 8'd59;8'd36: cx <= 8'd60;8'd37: cx <= 8'd60;8'd38: cx <= 8'd61;8'd39: cx <= 8'd62;8'd40: cx <= 8'd63;8'd41: cx <= 8'd63;8'd42: cx <= 8'd64;8'd43: cx <= 8'd65;8'd44: cx <= 8'd66;8'd45: cx <= 8'd66;8'd46: cx <= 8'd67;8'd47: cx <= 8'd68;8'd48: cx <= 8'd69;8'd49: cx <= 8'd69;8'd50: cx <= 8'd70;8'd51: cx <= 8'd71;8'd52: cx <= 8'd71;8'd53: cx <= 8'd72;8'd54: cx <= 8'd73;8'd55: cx <= 8'd74;8'd56: cx <= 8'd74;8'd57: cx <= 8'd75;8'd58: cx <= 8'd76;8'd59: cx <= 8'd77;8'd60: cx <= 8'd77;8'd61: cx <= 8'd78;8'd62: cx <= 8'd79;8'd63: cx <= 8'd80;8'd64: cx <= 8'd80;8'd65: cx <= 8'd81;8'd66: cx <= 8'd82;8'd67: cx <= 8'd83;8'd68: cx <= 8'd83;8'd69: cx <= 8'd84;8'd70: cx <= 8'd85;8'd71: cx <= 8'd86;8'd72: cx <= 8'd86;8'd73: cx <= 8'd87;8'd74: cx <= 8'd88;8'd75: cx <= 8'd89;8'd76: cx <= 8'd89;8'd77: cx <= 8'd90;8'd78: cx <= 8'd91;8'd79: cx <= 8'd91;8'd80: cx <= 8'd92;8'd81: cx <= 8'd93;8'd82: cx <= 8'd94;8'd83: cx <= 8'd94;8'd84: cx <= 8'd95;8'd85: cx <= 8'd96;8'd86: cx <= 8'd97;8'd87: cx <= 8'd97;8'd88: cx <= 8'd98;8'd89: cx <= 8'd99;8'd90: cx <= 8'd100;8'd91: cx <= 8'd100;8'd92: cx <= 8'd101;8'd93: cx <= 8'd102;8'd94: cx <= 8'd103;8'd95: cx <= 8'd103;8'd96: cx <= 8'd104;8'd97: cx <= 8'd105;8'd98: cx <= 8'd106;8'd99: cx <= 8'd106;8'd100: cx <= 8'd107;8'd101: cx <= 8'd108;8'd102: cx <= 8'd108;8'd103: cx <= 8'd109;8'd104: cx <= 8'd110;8'd105: cx <= 8'd111;8'd106: cx <= 8'd111;8'd107: cx <= 8'd112;8'd108: cx <= 8'd113;8'd109: cx <= 8'd114;8'd110: cx <= 8'd114;8'd111: cx <= 8'd115;8'd112: cx <= 8'd116;8'd113: cx <= 8'd117;8'd114: cx <= 8'd117;8'd115: cx <= 8'd118;8'd116: cx <= 8'd119;8'd117: cx <= 8'd120;8'd118: cx <= 8'd120;8'd119: cx <= 8'd121;8'd120: cx <= 8'd122;8'd121: cx <= 8'd123;8'd122: cx <= 8'd123;8'd123: cx <= 8'd124;8'd124: cx <= 8'd125;8'd125: cx <= 8'd126;8'd126: cx <= 8'd126;8'd127: cx <= 8'd127;8'd128: cx <= 8'd128;8'd129: cx <= 8'd128;8'd130: cx <= 8'd129;8'd131: cx <= 8'd130;8'd132: cx <= 8'd131;8'd133: cx <= 8'd131;8'd134: cx <= 8'd132;8'd135: cx <= 8'd133;8'd136: cx <= 8'd134;8'd137: cx <= 8'd134;8'd138: cx <= 8'd135;8'd139: cx <= 8'd136;8'd140: cx <= 8'd137;8'd141: cx <= 8'd137;8'd142: cx <= 8'd138;8'd143: cx <= 8'd139;8'd144: cx <= 8'd140;8'd145: cx <= 8'd140;8'd146: cx <= 8'd141;8'd147: cx <= 8'd142;8'd148: cx <= 8'd143;8'd149: cx <= 8'd143;8'd150: cx <= 8'd144;8'd151: cx <= 8'd145;8'd152: cx <= 8'd146;8'd153: cx <= 8'd146;8'd154: cx <= 8'd147;8'd155: cx <= 8'd148;8'd156: cx <= 8'd148;8'd157: cx <= 8'd149;8'd158: cx <= 8'd150;8'd159: cx <= 8'd151;8'd160: cx <= 8'd151;8'd161: cx <= 8'd152;8'd162: cx <= 8'd153;8'd163: cx <= 8'd154;8'd164: cx <= 8'd154;8'd165: cx <= 8'd155;8'd166: cx <= 8'd156;8'd167: cx <= 8'd157;8'd168: cx <= 8'd157;8'd169: cx <= 8'd158;8'd170: cx <= 8'd159;8'd171: cx <= 8'd160;8'd172: cx <= 8'd160;8'd173: cx <= 8'd161;8'd174: cx <= 8'd162;8'd175: cx <= 8'd163;8'd176: cx <= 8'd163;8'd177: cx <= 8'd164;8'd178: cx <= 8'd165;8'd179: cx <= 8'd165;8'd180: cx <= 8'd166;8'd181: cx <= 8'd167;8'd182: cx <= 8'd168;8'd183: cx <= 8'd168;8'd184: cx <= 8'd169;8'd185: cx <= 8'd170;8'd186: cx <= 8'd171;8'd187: cx <= 8'd171;8'd188: cx <= 8'd172;8'd189: cx <= 8'd173;8'd190: cx <= 8'd174;8'd191: cx <= 8'd174;8'd192: cx <= 8'd175;8'd193: cx <= 8'd176;8'd194: cx <= 8'd177;8'd195: cx <= 8'd177;8'd196: cx <= 8'd178;8'd197: cx <= 8'd179;8'd198: cx <= 8'd180;8'd199: cx <= 8'd180;8'd200: cx <= 8'd181;8'd201: cx <= 8'd182;8'd202: cx <= 8'd183;8'd203: cx <= 8'd183;8'd204: cx <= 8'd184;8'd205: cx <= 8'd185;8'd206: cx <= 8'd185;8'd207: cx <= 8'd186;8'd208: cx <= 8'd187;8'd209: cx <= 8'd188;8'd210: cx <= 8'd188;8'd211: cx <= 8'd189;8'd212: cx <= 8'd190;8'd213: cx <= 8'd191;8'd214: cx <= 8'd191;8'd215: cx <= 8'd192;8'd216: cx <= 8'd193;8'd217: cx <= 8'd194;8'd218: cx <= 8'd194;8'd219: cx <= 8'd195;8'd220: cx <= 8'd196;8'd221: cx <= 8'd197;8'd222: cx <= 8'd197;8'd223: cx <= 8'd198;8'd224: cx <= 8'd199;8'd225: cx <= 8'd200;8'd226: cx <= 8'd200;8'd227: cx <= 8'd201;8'd228: cx <= 8'd202;8'd229: cx <= 8'd202;8'd230: cx <= 8'd203;8'd231: cx <= 8'd204;8'd232: cx <= 8'd205;8'd233: cx <= 8'd205;8'd234: cx <= 8'd206;8'd235: cx <= 8'd207;8'd236: cx <= 8'd208;8'd237: cx <= 8'd208;8'd238: cx <= 8'd209;8'd239: cx <= 8'd210;8'd240: cx <= 8'd211;8'd241: cx <= 8'd211;8'd242: cx <= 8'd212;8'd243: cx <= 8'd213;8'd244: cx <= 8'd214;8'd245: cx <= 8'd214;8'd246: cx <= 8'd215;8'd247: cx <= 8'd216;8'd248: cx <= 8'd217;8'd249: cx <= 8'd217;8'd250: cx <= 8'd218;8'd251: cx <= 8'd219;8'd252: cx <= 8'd220;8'd253: cx <= 8'd220;8'd254: cx <= 8'd221;8'd255: cx <= 8'd222;default: cx<=8'd127; endcase case ( cycal )8'd0: cy <= 8'd33;8'd1: cy <= 8'd34;8'd2: cy <= 8'd34;8'd3: cy <= 8'd35;8'd4: cy <= 8'd36;8'd5: cy <= 8'd37;8'd6: cy <= 8'd37;8'd7: cy <= 8'd38;8'd8: cy <= 8'd39;8'd9: cy <= 8'd40;8'd10: cy <= 8'd40;8'd11: cy <= 8'd41;8'd12: cy <= 8'd42;8'd13: cy <= 8'd43;8'd14: cy <= 8'd43;8'd15: cy <= 8'd44;8'd16: cy <= 8'd45;8'd17: cy <= 8'd46;8'd18: cy <= 8'd46;8'd19: cy <= 8'd47;8'd20: cy <= 8'd48;8'd21: cy <= 8'd49;8'd22: cy <= 8'd49;8'd23: cy <= 8'd50;8'd24: cy <= 8'd51;8'd25: cy <= 8'd52;8'd26: cy <= 8'd52;8'd27: cy <= 8'd53;8'd28: cy <= 8'd54;8'd29: cy <= 8'd54;8'd30: cy <= 8'd55;8'd31: cy <= 8'd56;8'd32: cy <= 8'd57;8'd33: cy <= 8'd57;8'd34: cy <= 8'd58;8'd35: cy <= 8'd59;8'd36: cy <= 8'd60;8'd37: cy <= 8'd60;8'd38: cy <= 8'd61;8'd39: cy <= 8'd62;8'd40: cy <= 8'd63;8'd41: cy <= 8'd63;8'd42: cy <= 8'd64;8'd43: cy <= 8'd65;8'd44: cy <= 8'd66;8'd45: cy <= 8'd66;8'd46: cy <= 8'd67;8'd47: cy <= 8'd68;8'd48: cy <= 8'd69;8'd49: cy <= 8'd69;8'd50: cy <= 8'd70;8'd51: cy <= 8'd71;8'd52: cy <= 8'd71;8'd53: cy <= 8'd72;8'd54: cy <= 8'd73;8'd55: cy <= 8'd74;8'd56: cy <= 8'd74;8'd57: cy <= 8'd75;8'd58: cy <= 8'd76;8'd59: cy <= 8'd77;8'd60: cy <= 8'd77;8'd61: cy <= 8'd78;8'd62: cy <= 8'd79;8'd63: cy <= 8'd80;8'd64: cy <= 8'd80;8'd65: cy <= 8'd81;8'd66: cy <= 8'd82;8'd67: cy <= 8'd83;8'd68: cy <= 8'd83;8'd69: cy <= 8'd84;8'd70: cy <= 8'd85;8'd71: cy <= 8'd86;8'd72: cy <= 8'd86;8'd73: cy <= 8'd87;8'd74: cy <= 8'd88;8'd75: cy <= 8'd89;8'd76: cy <= 8'd89;8'd77: cy <= 8'd90;8'd78: cy <= 8'd91;8'd79: cy <= 8'd91;8'd80: cy <= 8'd92;8'd81: cy <= 8'd93;8'd82: cy <= 8'd94;8'd83: cy <= 8'd94;8'd84: cy <= 8'd95;8'd85: cy <= 8'd96;8'd86: cy <= 8'd97;8'd87: cy <= 8'd97;8'd88: cy <= 8'd98;8'd89: cy <= 8'd99;8'd90: cy <= 8'd100;8'd91: cy <= 8'd100;8'd92: cy <= 8'd101;8'd93: cy <= 8'd102;8'd94: cy <= 8'd103;8'd95: cy <= 8'd103;8'd96: cy <= 8'd104;8'd97: cy <= 8'd105;8'd98: cy <= 8'd106;8'd99: cy <= 8'd106;8'd100: cy <= 8'd107;8'd101: cy <= 8'd108;8'd102: cy <= 8'd108;8'd103: cy <= 8'd109;8'd104: cy <= 8'd110;8'd105: cy <= 8'd111;8'd106: cy <= 8'd111;8'd107: cy <= 8'd112;8'd108: cy <= 8'd113;8'd109: cy <= 8'd114;8'd110: cy <= 8'd114;8'd111: cy <= 8'd115;8'd112: cy <= 8'd116;8'd113: cy <= 8'd117;8'd114: cy <= 8'd117;8'd115: cy <= 8'd118;8'd116: cy <= 8'd119;8'd117: cy <= 8'd120;8'd118: cy <= 8'd120;8'd119: cy <= 8'd121;8'd120: cy <= 8'd122;8'd121: cy <= 8'd123;8'd122: cy <= 8'd123;8'd123: cy <= 8'd124;8'd124: cy <= 8'd125;8'd125: cy <= 8'd126;8'd126: cy <= 8'd126;8'd127: cy <= 8'd127;8'd128: cy <= 8'd128;8'd129: cy <= 8'd128;8'd130: cy <= 8'd129;8'd131: cy <= 8'd130;8'd132: cy <= 8'd131;8'd133: cy <= 8'd131;8'd134: cy <= 8'd132;8'd135: cy <= 8'd133;8'd136: cy <= 8'd134;8'd137: cy <= 8'd134;8'd138: cy <= 8'd135;8'd139: cy <= 8'd136;8'd140: cy <= 8'd137;8'd141: cy <= 8'd137;8'd142: cy <= 8'd138;8'd143: cy <= 8'd139;8'd144: cy <= 8'd140;8'd145: cy <= 8'd140;8'd146: cy <= 8'd141;8'd147: cy <= 8'd142;8'd148: cy <= 8'd143;8'd149: cy <= 8'd143;8'd150: cy <= 8'd144;8'd151: cy <= 8'd145;8'd152: cy <= 8'd146;8'd153: cy <= 8'd146;8'd154: cy <= 8'd147;8'd155: cy <= 8'd148;8'd156: cy <= 8'd148;8'd157: cy <= 8'd149;8'd158: cy <= 8'd150;8'd159: cy <= 8'd151;8'd160: cy <= 8'd151;8'd161: cy <= 8'd152;8'd162: cy <= 8'd153;8'd163: cy <= 8'd154;8'd164: cy <= 8'd154;8'd165: cy <= 8'd155;8'd166: cy <= 8'd156;8'd167: cy <= 8'd157;8'd168: cy <= 8'd157;8'd169: cy <= 8'd158;8'd170: cy <= 8'd159;8'd171: cy <= 8'd160;8'd172: cy <= 8'd160;8'd173: cy <= 8'd161;8'd174: cy <= 8'd162;8'd175: cy <= 8'd163;8'd176: cy <= 8'd163;8'd177: cy <= 8'd164;8'd178: cy <= 8'd165;8'd179: cy <= 8'd165;8'd180: cy <= 8'd166;8'd181: cy <= 8'd167;8'd182: cy <= 8'd168;8'd183: cy <= 8'd168;8'd184: cy <= 8'd169;8'd185: cy <= 8'd170;8'd186: cy <= 8'd171;8'd187: cy <= 8'd171;8'd188: cy <= 8'd172;8'd189: cy <= 8'd173;8'd190: cy <= 8'd174;8'd191: cy <= 8'd174;8'd192: cy <= 8'd175;8'd193: cy <= 8'd176;8'd194: cy <= 8'd177;8'd195: cy <= 8'd177;8'd196: cy <= 8'd178;8'd197: cy <= 8'd179;8'd198: cy <= 8'd180;8'd199: cy <= 8'd180;8'd200: cy <= 8'd181;8'd201: cy <= 8'd182;8'd202: cy <= 8'd183;8'd203: cy <= 8'd183;8'd204: cy <= 8'd184;8'd205: cy <= 8'd185;8'd206: cy <= 8'd185;8'd207: cy <= 8'd186;8'd208: cy <= 8'd187;8'd209: cy <= 8'd188;8'd210: cy <= 8'd188;8'd211: cy <= 8'd189;8'd212: cy <= 8'd190;8'd213: cy <= 8'd191;8'd214: cy <= 8'd191;8'd215: cy <= 8'd192;8'd216: cy <= 8'd193;8'd217: cy <= 8'd194;8'd218: cy <= 8'd194;8'd219: cy <= 8'd195;8'd220: cy <= 8'd196;8'd221: cy <= 8'd197;8'd222: cy <= 8'd197;8'd223: cy <= 8'd198;8'd224: cy <= 8'd199;8'd225: cy <= 8'd200;8'd226: cy <= 8'd200;8'd227: cy <= 8'd201;8'd228: cy <= 8'd202;8'd229: cy <= 8'd202;8'd230: cy <= 8'd203;8'd231: cy <= 8'd204;8'd232: cy <= 8'd205;8'd233: cy <= 8'd205;8'd234: cy <= 8'd206;8'd235: cy <= 8'd207;8'd236: cy <= 8'd208;8'd237: cy <= 8'd208;8'd238: cy <= 8'd209;8'd239: cy <= 8'd210;8'd240: cy <= 8'd211;8'd241: cy <= 8'd211;8'd242: cy <= 8'd212;8'd243: cy <= 8'd213;8'd244: cy <= 8'd214;8'd245: cy <= 8'd214;8'd246: cy <= 8'd215;8'd247: cy <= 8'd216;8'd248: cy <= 8'd217;8'd249: cy <= 8'd217;8'd250: cy <= 8'd218;8'd251: cy <= 8'd219;8'd252: cy <= 8'd220;8'd253: cy <= 8'd220;8'd254: cy <= 8'd221;8'd255: cy <= 8'd222;default: cy<=8'd127; endcase 

    if ( connected == 1 ) begin
        GCBD[15:0] <= GCdata[64:49]; //button data
        if ( NSOCal == 0 ) begin // 0 is when button is held to enter NSO MODE
            GCLA[15:0] <= {  x[7:0] , y[7:0]  };
            GCRA[15:0] <= { cx[7:0] , cy[7:0] };
        end else begin
            GCLA[15:0] <= {  xcal[7:0] , ycal[7:0] };   //GCdata[48:41] , GCdata[40:33] };          //{ $signed({1'b0,GCdata[48:41]})-$signed(offsetx) , $signed({1'b0,GCdata[40:33]})-$signed(offsety) };
            GCRA[15:0] <= { cxcal[7:0] ,cycal[7:0] };   //GCdata[32:25] , GCdata[24:17] };          //{ $signed({1'b0,GCdata[32:25]})-$signed(offsetcx) , $signed({1'b0,GCdata[24:17]})-$signed(offsetcy) }; 
        end
    end
    else begin
        GCBD[15:0] <= 16'h0000;
        x[7:0] <= 8'h7F;
        y[7:0] <= 8'h7F;
        cx[7:0]<= 8'h7F;
        cy[7:0]<= 8'h7F;
    end
    if ( ( {1'b0,GCdata[16:09]} - $signed(offsetLT) ) > 8'b11111111 ) begin
        LAT[7:0] <= 8'b0;
    end else begin
        LAT[7:0] <= GCdata[16:09] - $signed(offsetLT);
    end
    if ( ( {1'b0,GCdata[08:01]} - $signed(offsetRT) ) > 8'b11111111 ) begin
        RAT[7:0] <= 8'b0;
    end else begin
        RAT[7:0] <= GCdata[08:01] - $signed(offsetRT);
    end
    GCTA[15:0] = {LAT[7:0] , RAT[7:0]};
end

reg [81:0] GCdata = 82'b0;
always @ ( posedge clk ) begin

    prev_POLL <= POLL;

    if ( GC_enable == 1 ) begin

        if ( prev_POLL && ~POLL ) begin // falling edge detected
            count <= 1'b0;
            bit_count <= bit_count - 1'b1;
        end

        if ( ~prev_POLL && ~POLL ) begin // controller line low
            count <= count + 1'b1;
        end

        if ( ~prev_POLL && POLL ) begin // rising edge detected
            if ( count > 55 ) begin              
                GCdata[81:0] <= (GCdata[81:0] << 1) | 1'b0 ;
                count <= 1'b0;
            end
            else begin
                GCdata[81:0] <= (GCdata[81:0] << 1) | 1'b1 ;
                count <= 1'b0;
            end
        end

        if ( prev_POLL && POLL ) begin // controller line high
            if ( count > 750 ) begin //F*** the Phob and ProGCC controllers. The delay to respond to the GC polling is so long it resets my counter. The delay is up to 24us. Fix your shit!
                GCpollend <= 1;
                if ( bit_count > 78 ) begin
                    connected <= 0;
                    connection_type <= 3'b000;
                end
                else if ( bit_count == 1 )begin
                    connected <= 0;
                    connection_type <= 3'b010;
                    NSOCal   <= button2;
                    offsetx  <= $signed({1'b0,GCdata[64:57]}) - 9'sd127;
                    offsety  <= $signed({1'b0,GCdata[56:49]}) - 9'sd127;
                    offsetcx <= $signed({1'b0,GCdata[48:41]}) - 9'sd127;
                    offsetcy <= $signed({1'b0,GCdata[40:33]}) - 9'sd127;
                    offsetLT <= GCdata[32:25];
                    offsetRT <= GCdata[24:17];
                end
                else if ( bit_count == 57 ) begin
                    connected <= 0;
                    connection_type <= 3'b001;
                end
                else if ( bit_count == 17 ) begin 
                    connected <= 1;
                    connection_type <= 3'b010;
                end
                else begin
                    connected <= 0;
                    connection_type <= 3'b000;
                end
            end
            else begin
                count <= count + 1'b1;
                GCpollend <= 0;
            end

        end

    end

    else begin  // if GC_enable is 0 then it is not the controller's turn to send data
        count <= 1'b0;
        prev_POLL <= 0; 
        bit_count <= 82;
    end
        
end
    

endmodule
